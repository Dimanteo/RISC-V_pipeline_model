module rv32(input clk, reset,
            output [31:0] pc,
            input [31:0] fetchI,
            output memWE,
            output [31:0] aluout, writedata,
            input [31:0] readdata);
    wire memtoreg, branch, alusrc, regdst, regwrite, writesmem,
         indirectbr, jump, invcond, uncond, genupimm, pcrel, pauseD;
    wire [3:0] alucontrol;
    wire [2:0] itype;
    wire [31:0] simm, uimm, decodeI;
    maindec md (.op(decodeI[6:0]),
                .funct3(decodeI[14:12]),
                .funct7(decodeI[31:25]),
                .memtoreg(memtoreg),
                .memwrite(writesmem),
                .alusrcimm(alusrc),
                .writesreg(regwrite),
                .indirectbr(indirectbr),
                .jump(jump),
                .pause(pauseD),
                .aluop(alucontrol), 
                .itype(itype),
                .invcond(invcond),
                .uncond(uncond),
                .genupimm(genupimm),
                .pcrel(pcrel));
    immdec immd(.instr(decodeI), .itype(itype), .simm(simm), .uimm(uimm));
    datapath dp(.clk(clk), .reset(reset), 
                .memtoreg(memtoreg),
                .alusrcimm(alusrc), 
                .writesreg(regwrite),
                .writesmem(writesmem),
                .indirectbr(indirectbr),
                .jump(jump),
                .invcond(invcond),
                .uncond(uncond),
                .genupimm(genupimm),
                .pcrel(pcrel),
                .pauseD(pauseD),
                .memWE(memWE),
                .simm(simm),
                .uimm(uimm),
                .alucontrol(alucontrol),
                .pc(pc), 
                .instr(fetchI),
                .decodeI(decodeI),
                .aluout(aluout),
                .writedata(writedata),
                .readdata(readdata));
endmodule