module adder(input [31:0] l, input [31:0] r, output [31:0] y);
    assign y = l + r;
endmodule